std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(129, 8)),
std_logic_vector(to_unsigned(130, 8)),
std_logic_vector(to_unsigned(132, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(135, 8)),
std_logic_vector(to_unsigned(136, 8)),
std_logic_vector(to_unsigned(138, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(141, 8)),
std_logic_vector(to_unsigned(143, 8)),
std_logic_vector(to_unsigned(144, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(147, 8)),
std_logic_vector(to_unsigned(149, 8)),
std_logic_vector(to_unsigned(150, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(153, 8)),
std_logic_vector(to_unsigned(155, 8)),
std_logic_vector(to_unsigned(156, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(159, 8)),
std_logic_vector(to_unsigned(161, 8)),
std_logic_vector(to_unsigned(162, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(165, 8)),
std_logic_vector(to_unsigned(167, 8)),
std_logic_vector(to_unsigned(168, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(171, 8)),
std_logic_vector(to_unsigned(173, 8)),
std_logic_vector(to_unsigned(174, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(177, 8)),
std_logic_vector(to_unsigned(178, 8)),
std_logic_vector(to_unsigned(180, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(183, 8)),
std_logic_vector(to_unsigned(184, 8)),
std_logic_vector(to_unsigned(185, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(188, 8)),
std_logic_vector(to_unsigned(190, 8)),
std_logic_vector(to_unsigned(191, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(194, 8)),
std_logic_vector(to_unsigned(195, 8)),
std_logic_vector(to_unsigned(196, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(199, 8)),
std_logic_vector(to_unsigned(200, 8)),
std_logic_vector(to_unsigned(201, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(204, 8)),
std_logic_vector(to_unsigned(205, 8)),
std_logic_vector(to_unsigned(206, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(209, 8)),
std_logic_vector(to_unsigned(210, 8)),
std_logic_vector(to_unsigned(211, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(213, 8)),
std_logic_vector(to_unsigned(215, 8)),
std_logic_vector(to_unsigned(216, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(218, 8)),
std_logic_vector(to_unsigned(219, 8)),
std_logic_vector(to_unsigned(220, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(222, 8)),
std_logic_vector(to_unsigned(223, 8)),
std_logic_vector(to_unsigned(224, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(226, 8)),
std_logic_vector(to_unsigned(227, 8)),
std_logic_vector(to_unsigned(228, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(230, 8)),
std_logic_vector(to_unsigned(231, 8)),
std_logic_vector(to_unsigned(232, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(234, 8)),
std_logic_vector(to_unsigned(235, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(237, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(241, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(243, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(246, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(246, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(243, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(241, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(237, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(235, 8)),
std_logic_vector(to_unsigned(234, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(232, 8)),
std_logic_vector(to_unsigned(231, 8)),
std_logic_vector(to_unsigned(230, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(228, 8)),
std_logic_vector(to_unsigned(227, 8)),
std_logic_vector(to_unsigned(226, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(224, 8)),
std_logic_vector(to_unsigned(223, 8)),
std_logic_vector(to_unsigned(222, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(220, 8)),
std_logic_vector(to_unsigned(219, 8)),
std_logic_vector(to_unsigned(218, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(216, 8)),
std_logic_vector(to_unsigned(215, 8)),
std_logic_vector(to_unsigned(213, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(211, 8)),
std_logic_vector(to_unsigned(210, 8)),
std_logic_vector(to_unsigned(209, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(206, 8)),
std_logic_vector(to_unsigned(205, 8)),
std_logic_vector(to_unsigned(204, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(201, 8)),
std_logic_vector(to_unsigned(200, 8)),
std_logic_vector(to_unsigned(199, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(196, 8)),
std_logic_vector(to_unsigned(195, 8)),
std_logic_vector(to_unsigned(194, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(191, 8)),
std_logic_vector(to_unsigned(190, 8)),
std_logic_vector(to_unsigned(188, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(185, 8)),
std_logic_vector(to_unsigned(184, 8)),
std_logic_vector(to_unsigned(183, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(180, 8)),
std_logic_vector(to_unsigned(178, 8)),
std_logic_vector(to_unsigned(177, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(174, 8)),
std_logic_vector(to_unsigned(173, 8)),
std_logic_vector(to_unsigned(171, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(168, 8)),
std_logic_vector(to_unsigned(167, 8)),
std_logic_vector(to_unsigned(165, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(162, 8)),
std_logic_vector(to_unsigned(161, 8)),
std_logic_vector(to_unsigned(159, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(156, 8)),
std_logic_vector(to_unsigned(155, 8)),
std_logic_vector(to_unsigned(153, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(150, 8)),
std_logic_vector(to_unsigned(149, 8)),
std_logic_vector(to_unsigned(147, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(144, 8)),
std_logic_vector(to_unsigned(143, 8)),
std_logic_vector(to_unsigned(141, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(138, 8)),
std_logic_vector(to_unsigned(136, 8)),
std_logic_vector(to_unsigned(135, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(132, 8)),
std_logic_vector(to_unsigned(130, 8)),
std_logic_vector(to_unsigned(129, 8)),
std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(125, 8)),
std_logic_vector(to_unsigned(124, 8)),
std_logic_vector(to_unsigned(122, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(119, 8)),
std_logic_vector(to_unsigned(118, 8)),
std_logic_vector(to_unsigned(116, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(113, 8)),
std_logic_vector(to_unsigned(111, 8)),
std_logic_vector(to_unsigned(110, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(107, 8)),
std_logic_vector(to_unsigned(105, 8)),
std_logic_vector(to_unsigned(104, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(101, 8)),
std_logic_vector(to_unsigned(99, 8)),
std_logic_vector(to_unsigned(98, 8)),
std_logic_vector(to_unsigned(96, 8)),
std_logic_vector(to_unsigned(95, 8)),
std_logic_vector(to_unsigned(93, 8)),
std_logic_vector(to_unsigned(92, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(89, 8)),
std_logic_vector(to_unsigned(87, 8)),
std_logic_vector(to_unsigned(86, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(83, 8)),
std_logic_vector(to_unsigned(81, 8)),
std_logic_vector(to_unsigned(80, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(77, 8)),
std_logic_vector(to_unsigned(76, 8)),
std_logic_vector(to_unsigned(74, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(71, 8)),
std_logic_vector(to_unsigned(70, 8)),
std_logic_vector(to_unsigned(69, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(66, 8)),
std_logic_vector(to_unsigned(64, 8)),
std_logic_vector(to_unsigned(63, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(60, 8)),
std_logic_vector(to_unsigned(59, 8)),
std_logic_vector(to_unsigned(58, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(55, 8)),
std_logic_vector(to_unsigned(54, 8)),
std_logic_vector(to_unsigned(53, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(50, 8)),
std_logic_vector(to_unsigned(49, 8)),
std_logic_vector(to_unsigned(48, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(45, 8)),
std_logic_vector(to_unsigned(44, 8)),
std_logic_vector(to_unsigned(43, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(41, 8)),
std_logic_vector(to_unsigned(39, 8)),
std_logic_vector(to_unsigned(38, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(36, 8)),
std_logic_vector(to_unsigned(35, 8)),
std_logic_vector(to_unsigned(34, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(32, 8)),
std_logic_vector(to_unsigned(31, 8)),
std_logic_vector(to_unsigned(30, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(28, 8)),
std_logic_vector(to_unsigned(27, 8)),
std_logic_vector(to_unsigned(26, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(24, 8)),
std_logic_vector(to_unsigned(23, 8)),
std_logic_vector(to_unsigned(22, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(20, 8)),
std_logic_vector(to_unsigned(19, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(17, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(13, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(11, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(8, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(8, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(11, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(13, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(17, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(19, 8)),
std_logic_vector(to_unsigned(20, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(22, 8)),
std_logic_vector(to_unsigned(23, 8)),
std_logic_vector(to_unsigned(24, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(26, 8)),
std_logic_vector(to_unsigned(27, 8)),
std_logic_vector(to_unsigned(28, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(30, 8)),
std_logic_vector(to_unsigned(31, 8)),
std_logic_vector(to_unsigned(32, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(34, 8)),
std_logic_vector(to_unsigned(35, 8)),
std_logic_vector(to_unsigned(36, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(38, 8)),
std_logic_vector(to_unsigned(39, 8)),
std_logic_vector(to_unsigned(41, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(43, 8)),
std_logic_vector(to_unsigned(44, 8)),
std_logic_vector(to_unsigned(45, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(48, 8)),
std_logic_vector(to_unsigned(49, 8)),
std_logic_vector(to_unsigned(50, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(53, 8)),
std_logic_vector(to_unsigned(54, 8)),
std_logic_vector(to_unsigned(55, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(58, 8)),
std_logic_vector(to_unsigned(59, 8)),
std_logic_vector(to_unsigned(60, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(63, 8)),
std_logic_vector(to_unsigned(64, 8)),
std_logic_vector(to_unsigned(66, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(69, 8)),
std_logic_vector(to_unsigned(70, 8)),
std_logic_vector(to_unsigned(71, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(74, 8)),
std_logic_vector(to_unsigned(76, 8)),
std_logic_vector(to_unsigned(77, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(80, 8)),
std_logic_vector(to_unsigned(81, 8)),
std_logic_vector(to_unsigned(83, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(86, 8)),
std_logic_vector(to_unsigned(87, 8)),
std_logic_vector(to_unsigned(89, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(92, 8)),
std_logic_vector(to_unsigned(93, 8)),
std_logic_vector(to_unsigned(95, 8)),
std_logic_vector(to_unsigned(96, 8)),
std_logic_vector(to_unsigned(98, 8)),
std_logic_vector(to_unsigned(99, 8)),
std_logic_vector(to_unsigned(101, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(104, 8)),
std_logic_vector(to_unsigned(105, 8)),
std_logic_vector(to_unsigned(107, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(110, 8)),
std_logic_vector(to_unsigned(111, 8)),
std_logic_vector(to_unsigned(113, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(116, 8)),
std_logic_vector(to_unsigned(118, 8)),
std_logic_vector(to_unsigned(119, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(122, 8)),
std_logic_vector(to_unsigned(124, 8)),
std_logic_vector(to_unsigned(125, 8)),
std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(129, 8)),
std_logic_vector(to_unsigned(130, 8)),
std_logic_vector(to_unsigned(132, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(135, 8)),
std_logic_vector(to_unsigned(136, 8)),
std_logic_vector(to_unsigned(138, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(141, 8)),
std_logic_vector(to_unsigned(143, 8)),
std_logic_vector(to_unsigned(144, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(147, 8)),
std_logic_vector(to_unsigned(149, 8)),
std_logic_vector(to_unsigned(150, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(153, 8)),
std_logic_vector(to_unsigned(155, 8)),
std_logic_vector(to_unsigned(156, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(159, 8)),
std_logic_vector(to_unsigned(161, 8)),
std_logic_vector(to_unsigned(162, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(165, 8)),
std_logic_vector(to_unsigned(167, 8)),
std_logic_vector(to_unsigned(168, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(171, 8)),
std_logic_vector(to_unsigned(173, 8)),
std_logic_vector(to_unsigned(174, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(177, 8)),
std_logic_vector(to_unsigned(178, 8)),
std_logic_vector(to_unsigned(180, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(183, 8)),
std_logic_vector(to_unsigned(184, 8)),
std_logic_vector(to_unsigned(185, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(188, 8)),
std_logic_vector(to_unsigned(190, 8)),
std_logic_vector(to_unsigned(191, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(194, 8)),
std_logic_vector(to_unsigned(195, 8)),
std_logic_vector(to_unsigned(196, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(199, 8)),
std_logic_vector(to_unsigned(200, 8)),
std_logic_vector(to_unsigned(201, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(204, 8)),
std_logic_vector(to_unsigned(205, 8)),
std_logic_vector(to_unsigned(206, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(209, 8)),
std_logic_vector(to_unsigned(210, 8)),
std_logic_vector(to_unsigned(211, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(213, 8)),
std_logic_vector(to_unsigned(215, 8)),
std_logic_vector(to_unsigned(216, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(218, 8)),
std_logic_vector(to_unsigned(219, 8)),
std_logic_vector(to_unsigned(220, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(222, 8)),
std_logic_vector(to_unsigned(223, 8)),
std_logic_vector(to_unsigned(224, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(226, 8)),
std_logic_vector(to_unsigned(227, 8)),
std_logic_vector(to_unsigned(228, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(230, 8)),
std_logic_vector(to_unsigned(231, 8)),
std_logic_vector(to_unsigned(232, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(234, 8)),
std_logic_vector(to_unsigned(235, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(237, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(241, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(243, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(246, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(251, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(248, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(246, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(245, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(243, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(241, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(240, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(238, 8)),
std_logic_vector(to_unsigned(237, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(235, 8)),
std_logic_vector(to_unsigned(234, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(232, 8)),
std_logic_vector(to_unsigned(231, 8)),
std_logic_vector(to_unsigned(230, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(228, 8)),
std_logic_vector(to_unsigned(227, 8)),
std_logic_vector(to_unsigned(226, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(224, 8)),
std_logic_vector(to_unsigned(223, 8)),
std_logic_vector(to_unsigned(222, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(220, 8)),
std_logic_vector(to_unsigned(219, 8)),
std_logic_vector(to_unsigned(218, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(216, 8)),
std_logic_vector(to_unsigned(215, 8)),
std_logic_vector(to_unsigned(213, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(211, 8)),
std_logic_vector(to_unsigned(210, 8)),
std_logic_vector(to_unsigned(209, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(206, 8)),
std_logic_vector(to_unsigned(205, 8)),
std_logic_vector(to_unsigned(204, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(201, 8)),
std_logic_vector(to_unsigned(200, 8)),
std_logic_vector(to_unsigned(199, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(196, 8)),
std_logic_vector(to_unsigned(195, 8)),
std_logic_vector(to_unsigned(194, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(191, 8)),
std_logic_vector(to_unsigned(190, 8)),
std_logic_vector(to_unsigned(188, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(185, 8)),
std_logic_vector(to_unsigned(184, 8)),
std_logic_vector(to_unsigned(183, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(180, 8)),
std_logic_vector(to_unsigned(178, 8)),
std_logic_vector(to_unsigned(177, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(174, 8)),
std_logic_vector(to_unsigned(173, 8)),
std_logic_vector(to_unsigned(171, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(168, 8)),
std_logic_vector(to_unsigned(167, 8)),
std_logic_vector(to_unsigned(165, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(162, 8)),
std_logic_vector(to_unsigned(161, 8)),
std_logic_vector(to_unsigned(159, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(156, 8)),
std_logic_vector(to_unsigned(155, 8)),
std_logic_vector(to_unsigned(153, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(150, 8)),
std_logic_vector(to_unsigned(149, 8)),
std_logic_vector(to_unsigned(147, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(144, 8)),
std_logic_vector(to_unsigned(143, 8)),
std_logic_vector(to_unsigned(141, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(138, 8)),
std_logic_vector(to_unsigned(136, 8)),
std_logic_vector(to_unsigned(135, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(132, 8)),
std_logic_vector(to_unsigned(130, 8)),
std_logic_vector(to_unsigned(129, 8)),
std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(125, 8)),
std_logic_vector(to_unsigned(124, 8)),
std_logic_vector(to_unsigned(122, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(119, 8)),
std_logic_vector(to_unsigned(118, 8)),
std_logic_vector(to_unsigned(116, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(113, 8)),
std_logic_vector(to_unsigned(111, 8)),
std_logic_vector(to_unsigned(110, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(107, 8)),
std_logic_vector(to_unsigned(105, 8)),
std_logic_vector(to_unsigned(104, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(101, 8)),
std_logic_vector(to_unsigned(99, 8)),
std_logic_vector(to_unsigned(98, 8)),
std_logic_vector(to_unsigned(96, 8)),
std_logic_vector(to_unsigned(95, 8)),
std_logic_vector(to_unsigned(93, 8)),
std_logic_vector(to_unsigned(92, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(89, 8)),
std_logic_vector(to_unsigned(87, 8)),
std_logic_vector(to_unsigned(86, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(83, 8)),
std_logic_vector(to_unsigned(81, 8)),
std_logic_vector(to_unsigned(80, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(77, 8)),
std_logic_vector(to_unsigned(76, 8)),
std_logic_vector(to_unsigned(74, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(71, 8)),
std_logic_vector(to_unsigned(70, 8)),
std_logic_vector(to_unsigned(69, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(66, 8)),
std_logic_vector(to_unsigned(64, 8)),
std_logic_vector(to_unsigned(63, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(60, 8)),
std_logic_vector(to_unsigned(59, 8)),
std_logic_vector(to_unsigned(58, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(55, 8)),
std_logic_vector(to_unsigned(54, 8)),
std_logic_vector(to_unsigned(53, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(50, 8)),
std_logic_vector(to_unsigned(49, 8)),
std_logic_vector(to_unsigned(48, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(45, 8)),
std_logic_vector(to_unsigned(44, 8)),
std_logic_vector(to_unsigned(43, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(41, 8)),
std_logic_vector(to_unsigned(39, 8)),
std_logic_vector(to_unsigned(38, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(36, 8)),
std_logic_vector(to_unsigned(35, 8)),
std_logic_vector(to_unsigned(34, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(32, 8)),
std_logic_vector(to_unsigned(31, 8)),
std_logic_vector(to_unsigned(30, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(28, 8)),
std_logic_vector(to_unsigned(27, 8)),
std_logic_vector(to_unsigned(26, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(24, 8)),
std_logic_vector(to_unsigned(23, 8)),
std_logic_vector(to_unsigned(22, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(20, 8)),
std_logic_vector(to_unsigned(19, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(17, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(13, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(11, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(8, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(3, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(6, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(8, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(9, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(11, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(13, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(14, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(16, 8)),
std_logic_vector(to_unsigned(17, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(19, 8)),
std_logic_vector(to_unsigned(20, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(22, 8)),
std_logic_vector(to_unsigned(23, 8)),
std_logic_vector(to_unsigned(24, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(26, 8)),
std_logic_vector(to_unsigned(27, 8)),
std_logic_vector(to_unsigned(28, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(30, 8)),
std_logic_vector(to_unsigned(31, 8)),
std_logic_vector(to_unsigned(32, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(34, 8)),
std_logic_vector(to_unsigned(35, 8)),
std_logic_vector(to_unsigned(36, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(38, 8)),
std_logic_vector(to_unsigned(39, 8)),
std_logic_vector(to_unsigned(41, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(43, 8)),
std_logic_vector(to_unsigned(44, 8)),
std_logic_vector(to_unsigned(45, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(48, 8)),
std_logic_vector(to_unsigned(49, 8)),
std_logic_vector(to_unsigned(50, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(53, 8)),
std_logic_vector(to_unsigned(54, 8)),
std_logic_vector(to_unsigned(55, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(58, 8)),
std_logic_vector(to_unsigned(59, 8)),
std_logic_vector(to_unsigned(60, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(63, 8)),
std_logic_vector(to_unsigned(64, 8)),
std_logic_vector(to_unsigned(66, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(69, 8)),
std_logic_vector(to_unsigned(70, 8)),
std_logic_vector(to_unsigned(71, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(74, 8)),
std_logic_vector(to_unsigned(76, 8)),
std_logic_vector(to_unsigned(77, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(80, 8)),
std_logic_vector(to_unsigned(81, 8)),
std_logic_vector(to_unsigned(83, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(86, 8)),
std_logic_vector(to_unsigned(87, 8)),
std_logic_vector(to_unsigned(89, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(92, 8)),
std_logic_vector(to_unsigned(93, 8)),
std_logic_vector(to_unsigned(95, 8)),
std_logic_vector(to_unsigned(96, 8)),
std_logic_vector(to_unsigned(98, 8)),
std_logic_vector(to_unsigned(99, 8)),
std_logic_vector(to_unsigned(101, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(104, 8)),
std_logic_vector(to_unsigned(105, 8)),
std_logic_vector(to_unsigned(107, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(110, 8)),
std_logic_vector(to_unsigned(111, 8)),
std_logic_vector(to_unsigned(113, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(116, 8)),
std_logic_vector(to_unsigned(118, 8)),
std_logic_vector(to_unsigned(119, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(122, 8)),
std_logic_vector(to_unsigned(124, 8)),
std_logic_vector(to_unsigned(125, 8)),
